** Profile: "Ultrasonic_Generator-US_tran1"  [ D:\cad\cadence\EED3009-PSpiceFiles\Ultrasonic_Generator\US_tran1.sim ] 

** Creating circuit file "US_tran1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of D:\cad\cadence\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 50ms 0 1us 
.OPTIONS ADVCONV
.OPTIONS GMIN= 1.0E-9
.PROBE64 N([VOUT1])
.INC "..\Ultrasonic_Generator.net" 


.END
